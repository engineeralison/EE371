`timescale 1ns/1ps

module task2 (clk, reset, write, dataIn, address, dataOut);
	input logic clk, reset;
	input logic write;
	input logic [2:0] dataIn;
	input logic [4:0] address;
	output logic [2:0] dataOut;
	
	// 32x3 memory array
	logic [2:0] memory_array [31:0];
	
	logic [4:0] address_reg;
   logic [2:0] dataIn_reg;
   logic write_reg;
	
	// Register and pipeline the inputs
	always_ff @(posedge clk) begin
		if (reset) begin
			 address_reg <= 5'd0;
          dataIn_reg  <= 3'd0;
          write_reg   <= 1'b0;
        end 
        else begin
            address_reg <= address;
            dataIn_reg  <= dataIn;
            write_reg   <= write;
        end
    end
	 
	 // Write data into into memory array when write_reg is asserted
	  always_ff @(posedge clk) begin
        if (write_reg) begin
            memory_array[address_reg] <= dataIn_reg;
        end
    end
	 
	 // Read data out of the memory array
	 assign dataOut = memory_array[address_reg];
	
endmodule 