
module part2 (CLOCK_50, CLOCK2_50, KEY, SW, FPGA_I2C_SCLK, FPGA_I2C_SDAT, AUD_XCK, 
		        AUD_DACLRCK, AUD_ADCLRCK, AUD_BCLK, AUD_ADCDAT, AUD_DACDAT);

	// Clock signal inputs for system timing
	input CLOCK_50, CLOCK2_50;

	// Single-bit key input for reset functionality
	input [0:0] KEY;

	// 10-bit switch input for potential user interaction or control
	input [9:0] SW;

	// Audio/Video configuration interface using I2C protocol
	output FPGA_I2C_SCLK; // I2C clock signal
	inout FPGA_I2C_SDAT;  // I2C data signal

	// Audio codec interface signals
	output AUD_XCK;          // Audio clock signal
	input AUD_DACLRCK;       // DAC left/right clock
	input AUD_ADCLRCK;       // ADC left/right clock
	input AUD_BCLK;          // Audio bit clock
	input AUD_ADCDAT;        // ADC data input
	output AUD_DACDAT;       // DAC data output

	// Internal wires for handling read/write operations and data flow
	wire read_ready, write_ready;       // Flags for read/write readiness
	wire read, write;                   // Read and write control signals
	wire [23:0] readdata_left;          // Data read from the left audio channel
	wire [23:0] readdata_right;         // Data read from the right audio channel
	wire [23:0] writedata_left;         // Data to be written to the left audio channel
	wire [23:0] writedata_right;        // Data to be written to the right audio channel

	// Reset signal generated by inverting the key input
	wire reset = ~KEY[0];

	/////////////////////////////////
	// Your code goes here 
	/////////////////////////////////
	
	// Registers and wires for ROM data handling
	reg [15:0] rom_address;             // Address pointer for accessing ROM
	wire [23:0] data_from_rom;          // Data output from the ROM

	// Instantiation of the ROM module
	// ROM stores audio data that is read and processed for playback.
	note_data_ROM inst_ROM (
		.address(rom_address),          // Address input for ROM
		.clock(CLOCK_50),               // Clock input for synchronizing ROM operations
		.q(data_from_rom)               // Data output from ROM
	);

	// Sequential logic to manage ROM address updates
	always @(posedge CLOCK_50) begin
		 if (reset) begin
			rom_address <= 0;           // Reset the ROM address to the start
		 end
		 
		 if (write_ready) begin        // Update ROM address if write is ready
			  rom_address <= rom_address + 1; // Increment the ROM address
			  
			  if (rom_address >= 47_999) begin // Reset when reaching the max address
				rom_address <= 0;
			  end
		 end
	end

	// data to write to audio based off of switch condition
	assign writedata_left = SW[9] ? data_from_rom : readdata_left;
	assign writedata_right = SW[9] ? data_from_rom : readdata_right;
	
	// Write based off of switch 9 toggle
    assign write = SW[9] ? write_ready : (write_ready & read_ready);
	
	// Read based off of switch 9 toggle
    assign read = SW[9] ? read_ready : (write_ready & read_ready);
	
/////////////////////////////////////////////////////////////////////////////////
// Audio CODEC interface. 
//
// The interface consists of the following wires:
// read_ready, write_ready - CODEC ready for read/write operation 
// readdata_left, readdata_right - left and right channel data from the CODEC
// read - send data from the CODEC (both channels)
// writedata_left, writedata_right - left and right channel data to the CODEC
// write - send data to the CODEC (both channels)
// AUD_* - should connect to top-level entity I/O of the same name.
//         These signals go directly to the Audio CODEC
// I2C_* - should connect to top-level entity I/O of the same name.
//         These signals go directly to the Audio/Video Config module
/////////////////////////////////////////////////////////////////////////////////
	clock_generator my_clock_gen(
		// inputs
		CLOCK2_50,
		reset,

		// outputs
		AUD_XCK
	);

	audio_and_video_config cfg(
		// Inputs
		CLOCK_50,
		reset,

		// Bidirectionals
		FPGA_I2C_SDAT,
		FPGA_I2C_SCLK
	);

	audio_codec codec(
		// Inputs
		CLOCK_50,
		reset,

		read,	write,
		writedata_left, writedata_right,

		AUD_ADCDAT,

		// Bidirectionals
		AUD_BCLK,
		AUD_ADCLRCK,
		AUD_DACLRCK,

		// Outputs
		read_ready, write_ready,
		readdata_left, readdata_right,
		AUD_DACDAT
	);

endmodule